library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library math_library;
    use math_library.multiplier_pkg.all;

package field_oriented_motor_control_pkg is

end package field_oriented_motor_control_pkg;

package body field_oriented_motor_control_pkg is

end package body field_oriented_motor_control_pkg;
